// EMPTY !
// Need to specify directions and connections statically

module xmos_cpld_slice
(
// {ALTERA_ARGS_BEGIN} DO NOT REMOVE THIS LINE!

    AB10,
    AA11,
    AB11,
    AA12,
    AB12,
    AA13,
    CLK,
    AB13,
    AA15,
    AB15,
    AA16,
    AB17,
    nRST,
    B18,
    AA18,
    BA18,
    BB17,
    BA16,
    BB15,
    BA15,
    BB13,
    BA13,
    BB12,
    BA12,
    BB11,
    BA11,
    BB10,
    BA9,
    BB9,
    BA8,
    BB7,
    BA7,
    BB6,
    BA6,
    BB4,
    BA4,
    BB2,
    BA3,
    BB1,
    BA1,
    AA1,
    AB1,
    AA3,
    AB2,
    AA4,
    AB4,
    P55,
    AA6,
    AB6,
    AA7,
    AB7,
    AA8,
    AB9,
    AA9
// {ALTERA_ARGS_END} DO NOT REMOVE THIS LINE!

);

// {ALTERA_IO_BEGIN} DO NOT REMOVE THIS LINE!
inout           AB10;
inout           AA11;
inout           AB11;
inout           AA12;
inout           AB12;
inout           AA13;
input           CLK;
inout           AB13;
inout           AA15;
inout           AB15;
inout           AA16;
inout           AB17;
input           nRST;
input           B18;
inout           AA18;
inout           BA18;
inout           BB17;
inout           BA16;
inout           BB15;
inout           BA15;
inout           BB13;
inout           BA13;
inout           BB12;
inout           BA12;
inout           BB11;
inout           BA11;
input           BB10;
input           BA9;
input           BB9;
input           BA8;
input           BB7;
input           BA7;
input           BB6;
input           BA6;
input           BB4;
input           BA4;
input           BB2;
input           BA3;
input           BB1;
input           BA1;
input           AA1;
input           AB1;
input           AA3;
input           AB2;
input           AA4;
input           AB4;
input           P55;
input           AA6;
input           AB6;
input           AA7;
input           AB7;
inout           AA8;
input           AB9;
input           AA9;

// {ALTERA_IO_END} DO NOT REMOVE THIS LINE!
// {ALTERA_MODULE_BEGIN} DO NOT REMOVE THIS LINE!

// {ALTERA_MODULE_END} DO NOT REMOVE THIS LINE!
endmodule
